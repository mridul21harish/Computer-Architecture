`include "wallaceTreeMultiplier.v"

module top;

reg [31:0]A;
reg [31:0]B;
reg clk;
    
wire [63:0]C;

    	wallaceTreeMultiplier wtm(A, B, clk, C);
    	
    	always #5 clk = ~clk;

    	initial
    	begin
    	clk = 1'b0;

    	#5
        	A = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
        	B = 32'b0000_0000_0000_0000_0000_0000_0000_0100;
    	#100
    		$display("\t %d\t%d\t%d", A, B, C);
        	A = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
        	B = 32'b0000_0000_0000_0000_0000_0000_0100_0001;
    	#100
    		$display("\t %d\t%d\t%d", A, B, C);
        	A = 32'b0000_0000_0000_0000_0000_0000_1000_0000;
        	B = 32'b0000_0000_0000_0000_0000_0000_0000_0101;
    	#100
    		$display("\t %d\t%d\t%d", A, B, C);
        	A = 32'b0000_0000_0000_0000_0000_0010_0000_0011;
        	B = 32'b0000_0000_0000_0000_0000_0100_0000_1000;
    	#100
    		$display("\t %d\t%d\t%d", A, B, C);
        	A = 32'b0000_0000_0000_0000_0000_0000_0100_1001;
        	B = 32'b0000_0000_0000_0000_0000_0000_0001_0100;
        #100
        	$display("\t %d\t%d\t%d", A, B, C);
        #900
	$finish;
    	end

endmodule
